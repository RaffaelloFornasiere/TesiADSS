----------------------------------------------------------------------
entity randomcircuit is
	port (
		in0		: in  std_logic;
		in1		: in  std_logic;
		in2		: in  std_logic;
		in3		: in  std_logic;
		in4		: in  std_logic;
		in5		: in  std_logic;
		in6		: in  std_logic;
		out0		: out std_logic;
		out1		: out std_logic;
		out2		: out std_logic;
		out3		: out std_logic;
		out4		: out std_logic;
		out5		: out std_logic;
		out6		: out std_logic
	);
end randomcircuit;
----------------------------------------------------------------------

----------------------------------------------------------------------
architecture struct of randomcircuit is
	signal net_0		: std_logic;
	signal net_1		: std_logic;
	signal net_2		: std_logic;
	signal net_3		: std_logic;
	signal net_4		: std_logic;
	signal net_5		: std_logic;
	signal net_6		: std_logic;
	signal net_7		: std_logic;
	signal net_8		: std_logic;
	signal net_9		: std_logic;
	signal net_10		: std_logic;
	signal net_11		: std_logic;
	signal net_12		: std_logic;
	signal net_13		: std_logic;
	signal net_14		: std_logic;
	signal net_15		: std_logic;
	signal net_16		: std_logic;
	signal net_17		: std_logic;
	signal net_18		: std_logic;
	signal net_19		: std_logic;
	signal net_20		: std_logic;
	signal net_21		: std_logic;
	signal net_22		: std_logic;
	signal net_23		: std_logic;
	signal net_24		: std_logic;
	signal net_25		: std_logic;
	signal net_26		: std_logic;
	signal net_27		: std_logic;
	signal net_28		: std_logic;
	signal net_29		: std_logic;
	signal net_30		: std_logic;
	signal net_31		: std_logic;
	signal net_32		: std_logic;
	signal net_33		: std_logic;
	signal net_34		: std_logic;
	signal net_35		: std_logic;
	signal net_36		: std_logic;
	signal net_37		: std_logic;
	signal net_38		: std_logic;
	signal net_39		: std_logic;
	signal net_40		: std_logic;
	signal net_41		: std_logic;
	signal net_42		: std_logic;
	signal net_43		: std_logic;
	signal net_44		: std_logic;
	signal net_45		: std_logic;
	signal net_46		: std_logic;
	signal net_47		: std_logic;
begin
	net_41 <= in0;
	net_42 <= in1;
	net_43 <= in2;
	net_44 <= in3;
	net_45 <= in4;
	net_46 <= in5;
	net_47 <= in6;
	U36 : NOR4 port map(A1 => net_45, A2 => net_41, A3 => net_41, A4 => net_41, Z => net_34);
	U37 : NOT1 port map(A1 => net_43, Z => net_35);
	U38 : XOR3 port map(A1 => net_47, A2 => net_43, A3 => net_41, Z => net_36);
	U39 : XNOR2 port map(A1 => net_42, A2 => net_42, Z => net_37);
	U40 : XNOR2 port map(A1 => net_47, A2 => net_47, Z => net_38);
	U41 : OR2 port map(A1 => net_46, A2 => net_41, Z => net_39);
	U42 : NOT1 port map(A1 => net_44, Z => net_40);
	U27 : XNOR2 port map(A1 => net_38, A2 => net_47, Z => net_26);
	U28 : XOR3 port map(A1 => net_40, A2 => net_43, A3 => net_40, Z => net_27);
	U29 : OR3 port map(A1 => net_44, A2 => net_47, A3 => net_45, Z => net_28);
	U30 : AND2 port map(A1 => net_46, A2 => net_47, Z => net_29);
	U31 : AND4 port map(A1 => net_45, A2 => net_47, A3 => net_43, A4 => net_39, Z => net_30);
	U32 : AND2 port map(A1 => net_43, A2 => net_44, Z => net_31);
	U33 : NAND4 port map(A1 => net_34, A2 => net_44, A3 => net_42, A4 => net_37, Z => net_32);
	U34 : NAND4 port map(A1 => net_41, A2 => net_42, A3 => net_43, A4 => net_34, Z => net_33);
	U22 : OR2 port map(A1 => net_27, A2 => net_28, Z => net_21);
	U23 : NAND2 port map(A1 => net_33, A2 => net_44, Z => net_22);
	U24 : AND2 port map(A1 => net_43, A2 => net_35, Z => net_23);
	U25 : XNOR2 port map(A1 => net_26, A2 => net_38, Z => net_24);
	U26 : AND4 port map(A1 => net_30, A2 => net_46, A3 => net_40, A4 => net_39, Z => net_25);
	U17 : NOR4 port map(A1 => net_21, A2 => net_39, A3 => net_37, A4 => net_46, Z => net_16);
	U18 : XOR2 port map(A1 => net_34, A2 => net_35, Z => net_17);
	U19 : NOR4 port map(A1 => net_23, A2 => net_29, A3 => net_45, A4 => net_28, Z => net_18);
	U20 : XNOR2 port map(A1 => net_46, A2 => net_39, Z => net_19);
	U21 : NAND2 port map(A1 => net_36, A2 => net_38, Z => net_20);
	U12 : OR3 port map(A1 => net_42, A2 => net_38, A3 => net_18, Z => net_11);
	U13 : NOT1 port map(A1 => net_31, Z => net_12);
	U14 : XNOR2 port map(A1 => net_45, A2 => net_22, Z => net_13);
	U15 : NAND4 port map(A1 => net_18, A2 => net_46, A3 => net_24, A4 => net_20, Z => net_14);
	U16 : NOR2 port map(A1 => net_37, A2 => net_25, Z => net_15);
	U6 : XNOR2 port map(A1 => net_40, A2 => net_30, Z => net_5);
	U7 : NAND2 port map(A1 => net_14, A2 => net_16, Z => net_6);
	U8 : XOR2 port map(A1 => net_22, A2 => net_25, Z => net_7);
	U9 : NAND4 port map(A1 => net_15, A2 => net_24, A3 => net_32, A4 => net_36, Z => net_8);
	U10 : NOR3 port map(A1 => net_19, A2 => net_20, A3 => net_16, Z => net_9);
	U11 : NOR3 port map(A1 => net_16, A2 => net_17, A3 => net_17, Z => net_10);
	U1 : NOR4 port map(A1 => net_37, A2 => net_41, A3 => net_42, A4 => net_21, Z => net_0);
	U2 : XOR2 port map(A1 => net_5, A2 => net_12, Z => net_1);
	U3 : NOT1 port map(A1 => net_9, Z => net_2);
	U4 : XOR3 port map(A1 => net_7, A2 => net_8, A3 => net_10, Z => net_3);
	U5 : XOR2 port map(A1 => net_6, A2 => net_10, Z => net_4);
	out0 <= net_4;
	out1 <= net_1;
	out2 <= net_11;
	out3 <= net_13;
	out4 <= net_2;
	out5 <= net_3;
	out6 <= net_0;
end struct;
